`timescale 1ns / 1ps 
 module progmemory(clk, pc, inst); 
 	reg[27:0] pmemory[0:31]; output reg[27:0] inst; input wire[4:0]pc; input wire clk; initial begin 
pmemory[0]=28'b1110_00000000_00000100_00000000;
pmemory[1]=28'b1110_00000001_00000101_00000000;
pmemory[2]=28'b0001_00011111_00000001_00000000;
pmemory[3]=28'b1001_00000101_00011111_00000101;
pmemory[4]=28'b0001_00000111_00000000_00000000;
pmemory[5]=28'b0000_00000100_00001000_00000000;
pmemory[6]=28'b0000_00000100_00000110_00000000;
pmemory[7]=28'b1000_00000111_00001000_00000111;
pmemory[8]=28'b0001_00011111_00000001_00000000;
pmemory[9]=28'b1001_00000110_00011111_00000110;
pmemory[10]=28'b0110_00001011_00000111_00000000;
pmemory[11]=28'b0000_00000111_00001000_00000000;
pmemory[12]=28'b0001_00000111_00000000_00000000;
pmemory[13]=28'b0001_00011111_00000001_00000000;
pmemory[14]=28'b1001_00000101_00011111_00000101;
pmemory[15]=28'b0110_00010000_00000110_00000000;
pmemory[16]=28'b0010_00001000_00000101_00000000;
pmemory[17]=28'b1111_11111111_11111111_11111111;
end 
 		always @(*) begin 
 		inst = pmemory[pc]; end 
 endmodule 
